//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Wed Jan 30 16:11:33 2019
// Version: v11.9 SP2 11.9.2.1
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// simulate0
module simulate0(
    // Inputs
    CLKA,
    // Outputs
    data
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  CLKA;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output data;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   CLKA;
wire   data_net_0;
wire   myclock_0_GLA;
wire   myclock_0_LOCK;
wire   data_net_1;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire   VCC_net;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign VCC_net = 1'b1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign data_net_1 = data_net_0;
assign data       = data_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------myclock
myclock myclock_0(
        // Inputs
        .POWERDOWN ( VCC_net ),
        .CLKA      ( CLKA ),
        // Outputs
        .LOCK      ( myclock_0_LOCK ),
        .GLA       ( myclock_0_GLA ) 
        );

//--------test
test test_0(
        // Inputs
        .rst  ( myclock_0_LOCK ),
        .clk  ( myclock_0_GLA ),
        // Outputs
        .data ( data_net_0 ) 
        );


endmodule
